/*
  Author:Aniket Badhan
*/

program axiTestBench;

	axiEnv env;
	initial begin
		env = new();
		env.run();
	end

endprogram
